module fif_flush ();

endmodule
